--------------------------------------------------------------------------------
--             IntMultiplier_UsingDSP_24_24_48_unsigned_F400_uid4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_24_24_48_unsigned_F400_uid4 is
   port ( clk, rst, stall : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_24_24_48_unsigned_F400_uid4 is
signal XX_m5 :  std_logic_vector(23 downto 0);
signal YY_m5 :  std_logic_vector(23 downto 0);
signal DSP_bh6_ch0_0, DSP_bh6_ch0_0_d1 :  std_logic_vector(69 downto 0);
signal heap_bh6_w47_0 :  std_logic;
signal heap_bh6_w46_0 :  std_logic;
signal heap_bh6_w45_0 :  std_logic;
signal heap_bh6_w44_0 :  std_logic;
signal heap_bh6_w43_0 :  std_logic;
signal heap_bh6_w42_0 :  std_logic;
signal heap_bh6_w41_0 :  std_logic;
signal heap_bh6_w40_0 :  std_logic;
signal heap_bh6_w39_0 :  std_logic;
signal heap_bh6_w38_0 :  std_logic;
signal heap_bh6_w37_0 :  std_logic;
signal heap_bh6_w36_0 :  std_logic;
signal heap_bh6_w35_0 :  std_logic;
signal heap_bh6_w34_0 :  std_logic;
signal heap_bh6_w33_0 :  std_logic;
signal heap_bh6_w32_0 :  std_logic;
signal heap_bh6_w31_0 :  std_logic;
signal heap_bh6_w30_0 :  std_logic;
signal heap_bh6_w29_0 :  std_logic;
signal heap_bh6_w28_0 :  std_logic;
signal heap_bh6_w27_0 :  std_logic;
signal heap_bh6_w26_0 :  std_logic;
signal heap_bh6_w25_0 :  std_logic;
signal heap_bh6_w24_0 :  std_logic;
signal heap_bh6_w23_0 :  std_logic;
signal heap_bh6_w22_0 :  std_logic;
signal heap_bh6_w21_0 :  std_logic;
signal heap_bh6_w20_0 :  std_logic;
signal heap_bh6_w19_0 :  std_logic;
signal heap_bh6_w18_0 :  std_logic;
signal heap_bh6_w17_0 :  std_logic;
signal heap_bh6_w16_0 :  std_logic;
signal heap_bh6_w15_0 :  std_logic;
signal heap_bh6_w14_0 :  std_logic;
signal heap_bh6_w13_0 :  std_logic;
signal heap_bh6_w12_0 :  std_logic;
signal heap_bh6_w11_0 :  std_logic;
signal heap_bh6_w10_0 :  std_logic;
signal heap_bh6_w9_0 :  std_logic;
signal heap_bh6_w8_0 :  std_logic;
signal heap_bh6_w7_0 :  std_logic;
signal heap_bh6_w6_0 :  std_logic;
signal heap_bh6_w5_0 :  std_logic;
signal heap_bh6_w4_0 :  std_logic;
signal heap_bh6_w3_0 :  std_logic;
signal heap_bh6_w2_0 :  std_logic;
signal heap_bh6_w1_0 :  std_logic;
signal heap_bh6_w0_0 :  std_logic;
signal CompressionResult6 :  std_logic_vector(47 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then 
          if stall = '1' then
            DSP_bh6_ch0_0_d1 <=  DSP_bh6_ch0_0_d1;
          else 
            DSP_bh6_ch0_0_d1 <=  DSP_bh6_ch0_0;
          end if;
         end if;
      end process;
   XX_m5 <= X ;
   YY_m5 <= Y ;
   
   -- Beginning of code generated by BitHeap::generateCompressorVHDL
   -- code generated by BitHeap::generateSupertileVHDL()
   ----------------Synchro barrier, entering cycle 0----------------
   DSP_bh6_ch0_0 <= std_logic_vector(unsigned("" & XX_m5(23 downto 0) & "00000000000") * unsigned("" & YY_m5(23 downto 0) & "00000000000"));
   ----------------Synchro barrier, entering cycle 1----------------
   heap_bh6_w47_0 <= DSP_bh6_ch0_0_d1(69); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w46_0 <= DSP_bh6_ch0_0_d1(68); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w45_0 <= DSP_bh6_ch0_0_d1(67); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w44_0 <= DSP_bh6_ch0_0_d1(66); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w43_0 <= DSP_bh6_ch0_0_d1(65); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w42_0 <= DSP_bh6_ch0_0_d1(64); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w41_0 <= DSP_bh6_ch0_0_d1(63); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w40_0 <= DSP_bh6_ch0_0_d1(62); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w39_0 <= DSP_bh6_ch0_0_d1(61); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w38_0 <= DSP_bh6_ch0_0_d1(60); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w37_0 <= DSP_bh6_ch0_0_d1(59); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w36_0 <= DSP_bh6_ch0_0_d1(58); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w35_0 <= DSP_bh6_ch0_0_d1(57); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w34_0 <= DSP_bh6_ch0_0_d1(56); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w33_0 <= DSP_bh6_ch0_0_d1(55); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w32_0 <= DSP_bh6_ch0_0_d1(54); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w31_0 <= DSP_bh6_ch0_0_d1(53); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w30_0 <= DSP_bh6_ch0_0_d1(52); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w29_0 <= DSP_bh6_ch0_0_d1(51); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w28_0 <= DSP_bh6_ch0_0_d1(50); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w27_0 <= DSP_bh6_ch0_0_d1(49); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w26_0 <= DSP_bh6_ch0_0_d1(48); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w25_0 <= DSP_bh6_ch0_0_d1(47); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w24_0 <= DSP_bh6_ch0_0_d1(46); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w23_0 <= DSP_bh6_ch0_0_d1(45); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w22_0 <= DSP_bh6_ch0_0_d1(44); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w21_0 <= DSP_bh6_ch0_0_d1(43); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w20_0 <= DSP_bh6_ch0_0_d1(42); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w19_0 <= DSP_bh6_ch0_0_d1(41); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w18_0 <= DSP_bh6_ch0_0_d1(40); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w17_0 <= DSP_bh6_ch0_0_d1(39); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w16_0 <= DSP_bh6_ch0_0_d1(38); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w15_0 <= DSP_bh6_ch0_0_d1(37); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w14_0 <= DSP_bh6_ch0_0_d1(36); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w13_0 <= DSP_bh6_ch0_0_d1(35); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w12_0 <= DSP_bh6_ch0_0_d1(34); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w11_0 <= DSP_bh6_ch0_0_d1(33); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w10_0 <= DSP_bh6_ch0_0_d1(32); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w9_0 <= DSP_bh6_ch0_0_d1(31); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w8_0 <= DSP_bh6_ch0_0_d1(30); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w7_0 <= DSP_bh6_ch0_0_d1(29); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w6_0 <= DSP_bh6_ch0_0_d1(28); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w5_0 <= DSP_bh6_ch0_0_d1(27); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w4_0 <= DSP_bh6_ch0_0_d1(26); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w3_0 <= DSP_bh6_ch0_0_d1(25); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w2_0 <= DSP_bh6_ch0_0_d1(24); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w1_0 <= DSP_bh6_ch0_0_d1(23); -- cycle= 1 cp= 4.05e-10
   heap_bh6_w0_0 <= DSP_bh6_ch0_0_d1(22); -- cycle= 1 cp= 4.05e-10
   ----------------Synchro barrier, entering cycle 0----------------

   -- Adding the constant bits
      -- All the constant bits are zero, nothing to add

   ----------------Synchro barrier, entering cycle 1----------------
   CompressionResult6 <= heap_bh6_w47_0 & heap_bh6_w46_0 & heap_bh6_w45_0 & heap_bh6_w44_0 & heap_bh6_w43_0 & heap_bh6_w42_0 & heap_bh6_w41_0 & heap_bh6_w40_0 & heap_bh6_w39_0 & heap_bh6_w38_0 & heap_bh6_w37_0 & heap_bh6_w36_0 & heap_bh6_w35_0 & heap_bh6_w34_0 & heap_bh6_w33_0 & heap_bh6_w32_0 & heap_bh6_w31_0 & heap_bh6_w30_0 & heap_bh6_w29_0 & heap_bh6_w28_0 & heap_bh6_w27_0 & heap_bh6_w26_0 & heap_bh6_w25_0 & heap_bh6_w24_0 & heap_bh6_w23_0 & heap_bh6_w22_0 & heap_bh6_w21_0 & heap_bh6_w20_0 & heap_bh6_w19_0 & heap_bh6_w18_0 & heap_bh6_w17_0 & heap_bh6_w16_0 & heap_bh6_w15_0 & heap_bh6_w14_0 & heap_bh6_w13_0 & heap_bh6_w12_0 & heap_bh6_w11_0 & heap_bh6_w10_0 & heap_bh6_w9_0 & heap_bh6_w8_0 & heap_bh6_w7_0 & heap_bh6_w6_0 & heap_bh6_w5_0 & heap_bh6_w4_0 & heap_bh6_w3_0 & heap_bh6_w2_0 & heap_bh6_w1_0 & heap_bh6_w0_0;
   -- End of code generated by BitHeap::generateCompressorVHDL
   R <= CompressionResult6(47 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_33_f400_uid10
--                     (IntAdderClassical_33_F400_uid12)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_f400_uid10 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(32 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_f400_uid10 is
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   --Classical
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--                      FPMult_8_23_8_23_8_23_F400_uid2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2011
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMult_8_23_8_23_8_23_F400_uid2 is
   port ( clk, rst, stall : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FPMult_8_23_8_23_8_23_F400_uid2 is
   component IntMultiplier_UsingDSP_24_24_48_unsigned_F400_uid4 is
      port ( clk, rst, stall : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_f400_uid10 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(32 downto 0)   );
   end component;

signal sign, sign_d1, sign_d2 :  std_logic;
signal expX :  std_logic_vector(7 downto 0);
signal expY :  std_logic_vector(7 downto 0);
signal expSumPreSub :  std_logic_vector(9 downto 0);
signal bias :  std_logic_vector(9 downto 0);
signal expSum, expSum_d1 :  std_logic_vector(9 downto 0);
signal sigX :  std_logic_vector(23 downto 0);
signal sigY :  std_logic_vector(23 downto 0);
signal sigProd :  std_logic_vector(47 downto 0);
signal excSel :  std_logic_vector(3 downto 0);
signal exc, exc_d1, exc_d2 :  std_logic_vector(1 downto 0);
signal norm :  std_logic;
signal expPostNorm :  std_logic_vector(9 downto 0);
signal sigProdExt, sigProdExt_d1 :  std_logic_vector(47 downto 0);
signal expSig, expSig_d1 :  std_logic_vector(32 downto 0);
signal sticky, sticky_d1 :  std_logic;
signal guard :  std_logic;
signal round :  std_logic;
signal expSigPostRound :  std_logic_vector(32 downto 0);
signal excPostNorm :  std_logic_vector(1 downto 0);
signal finalExc :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then 
          if stall='1' then
            sign_d1       <= sign_d1      ;
            sign_d2       <= sign_d2      ;
            expSum_d1     <= expSum_d1    ;
            exc_d1        <= exc_d1       ;
            exc_d2        <= exc_d2       ;
            sigProdExt_d1 <= sigProdExt_d1;
            expSig_d1     <= expSig_d1    ;
            sticky_d1     <= sticky_d1    ;
          else 
            sign_d1 <=  sign;
            sign_d2 <=  sign_d1;
            expSum_d1 <=  expSum;
            exc_d1 <=  exc;
            exc_d2 <=  exc_d1;
            sigProdExt_d1 <=  sigProdExt;
            expSig_d1 <=  expSig;
            sticky_d1 <=  sticky;
           end if;
         end if;
      end process;
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   expSumPreSub <= ("00" & expX) + ("00" & expY);
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   expSum <= expSumPreSub - bias;
   ----------------Synchro barrier, entering cycle 0----------------
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_UsingDSP_24_24_48_unsigned_F400_uid4  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 stall=> stall,
                 R => sigProd,
                 X => sigX,
                 Y => sigY);
   ----------------Synchro barrier, entering cycle 1----------------
   ----------------Synchro barrier, entering cycle 0----------------
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel select 
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   ----------------Synchro barrier, entering cycle 1----------------
   norm <= sigProd(47);
   -- exponent update
   expPostNorm <= expSum_d1 + ("000000000" & norm);
   ----------------Synchro barrier, entering cycle 1----------------
   -- significand normalization shift
   sigProdExt <= sigProd(46 downto 0) & "0" when norm='1' else
                         sigProd(45 downto 0) & "00";
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24);
   ----------------Synchro barrier, entering cycle 2----------------
   guard <= '0' when sigProdExt_d1(23 downto 0)="000000000000000000000000" else '1';
   round <= sticky_d1 and ( (guard and not(sigProdExt_d1(25))) or (sigProdExt_d1(25) ))  ;
   RoundingAdder: IntAdder_33_f400_uid10  -- pipelineDepth=0 maxInDelay=8.43e-10
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => round,
                 R => expSigPostRound   ,
                 X => expSig_d1,
                 Y => "000000000000000000000000000000000");
   with expSigPostRound(32 downto 31) select
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_d2 select 
   finalExc <= exc_d2 when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign_d2 & expSigPostRound(30 downto 0);
end architecture;

