// =============================================================================
// Company      : University of Glasgow
// Author:        Waqar Nabi
// 
// Create Date  : 2014.12.04
// Design Name  : 
// Module Name  : counterSimple 
// Project Name : TyTra
// Target Devices: Stratix V (D5/D8) 
//
// Tool versions: 
// Dependencies : 
//
// Revision     : 
// Revision 0.01. File Created
// 
// =============================================================================

// =============================================================================
// General Description
// -----------------------------------------------------------------------------
// A general purpose N-bit wrap-around counter.
// synchronous reset
// 
//==============================================================================

module counterSimple
#(
// =============================================================================
// ** Parameters 
// =============================================================================
// Size of word (parent should over-write this if needeD)
  parameter N = 10 
)

(
// =============================================================================
// ** Ports 
// =============================================================================
  output reg  [N-1:0] y,
 
  input reset,
  input clk
);

// =============================================================================
// ** Procedures and assignments
// =============================================================================
always @(posedge clk)
  if (reset)
    y <= 0;
  else
    y <= y+1;

endmodule
